library verilog;
use verilog.vl_types.all;
entity noteIdentification is
    generic(
        Z               : integer := 0;
        C               : integer := 1;
        Cs              : integer := 2;
        D               : integer := 3;
        Ds              : integer := 4;
        E               : integer := 5;
        F               : integer := 6;
        Fs              : integer := 7;
        G               : integer := 8;
        Gs              : integer := 9;
        A               : integer := 10;
        As              : integer := 11;
        B               : integer := 12;
        Btwo            : integer := 42;
        GSfive          : integer := 283;
        DSfive          : integer := 212;
        Cthree          : integer := 44;
        Aone            : integer := 18;
        Ctwo            : integer := 22;
        Gthree          : integer := 66;
        CStwo           : integer := 23;
        Afive           : integer := 300;
        Cfour           : integer := 89;
        Bthree          : integer := 84;
        Gtwo            : integer := 33;
        AStwo           : integer := 39;
        FSone           : integer := 15;
        ASfour          : integer := 159;
        Afour           : integer := 150;
        Fone            : integer := 14;
        GSone           : integer := 17;
        Athree          : integer := 75;
        Done            : integer := 12;
        DSfour          : integer := 106;
        Dfive           : integer := 200;
        ASfive          : integer := 318;
        CSone           : integer := 11;
        CSfive          : integer := 189;
        Eone            : integer := 14;
        FSfive          : integer := 252;
        Gfive           : integer := 267;
        Cfive           : integer := 178;
        Atwo            : integer := 37;
        Efive           : integer := 225;
        Ffive           : integer := 238;
        Ftwo            : integer := 29;
        GStwo           : integer := 35;
        Bfive           : integer := 337;
        FSfour          : integer := 126;
        FSthree         : integer := 63;
        GSfour          : integer := 141;
        Ffour           : integer := 119;
        Dtwo            : integer := 25;
        Etwo            : integer := 28;
        Bfour           : integer := 168;
        DSone           : integer := 13;
        Ethree          : integer := 56;
        DStwo           : integer := 26;
        Fthree          : integer := 59;
        GSthree         : integer := 70;
        ASone           : integer := 19;
        FStwo           : integer := 31;
        Bone            : integer := 21;
        ASthree         : integer := 79;
        Gone            : integer := 16;
        CSfour          : integer := 94;
        Dfour           : integer := 100;
        Efour           : integer := 112;
        CSthree         : integer := 47;
        DSthree         : integer := 53;
        Gfour           : integer := 133;
        Cone            : integer := 11;
        Dthree          : integer := 50
    );
    port(
        reset           : in     vl_logic;
        clk             : in     vl_logic;
        ready           : in     vl_logic;
        switch          : in     vl_logic_vector(7 downto 0);
        from_ac97_data  : in     vl_logic_vector(15 downto 0);
        note            : out    vl_logic_vector(3 downto 0);
        GuessAddr       : out    vl_logic_vector(5 downto 0);
        readVal         : out    vl_logic;
        analyzer1_out   : out    vl_logic_vector(15 downto 0);
        analyzer2_out   : out    vl_logic_vector(15 downto 0)
    );
end noteIdentification;
